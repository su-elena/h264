`default_nettype none
`timescale 1ns / 1ps

module top_level(
    input wire clk,
    input wire btnc,
    output logic eth_rstn,
    output logic eth_txen,
    output wire eth_refclk, 
    output logic [1:0] eth_txd,
);

    
endmodule

`default nettype wire