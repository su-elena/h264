`default_nettype none
`timescale 1ns / 1ps

module chroma_subsample (
    input wire clk,
    input wire rst,
    input wire valid_in,
    input wire [19:0][14:0] addr,
    input wire [15:0][15:0] macroblock [23:0],
    output logic [15:0][15:0] macroblock_out [23:0],
    output logic [19:0][14:0] address,
    output wire valid_out
);
    logic [1:0][1:0][23:0] block1, block2, block3, block4, block5, block6, block7, block8;
    logic [1:0][15:0][23:0] row1;
    logic [1:0][1:0][23:0] block9, block10, block11, block12, block13, block14, block15, block16;
    logic [1:0][15:0][23:0] row2;
    logic [1:0][1:0][23:0] block17, block18, block19, block20, block21, block22, block23, block24;
    logic [1:0][15:0][23:0] row3;
    logic [1:0][1:0][23:0] block25, block26, block27, block28, block29, block30, block31, block32;
    logic [1:0][15:0][23:0] row4;
    logic [1:0][1:0][23:0] block33, block34, block35, block36, block37, block38, block39, block40;
    logic [1:0][15:0][23:0] row5;
    logic [1:0][1:0][23:0] block41, block42, block43, block44, block45, block46, block47, block48;
    logic [1:0][15:0][23:0] row6;
    logic [1:0][1:0][23:0] block49, block50, block51, block52, block53, block54, block55, block56;
    logic [1:0][15:0][23:0] row7;
    logic [1:0][1:0][23:0] block57, block58, block59, block60, block61, block62, block63, block64;
    logic [1:0][15:0][23:0] row8;

    logic prev_valid0, prev_valid1;

    always_ff @(posedge clk) begin
        prev_valid0 <= valid_in;
        prev_valid1 <= prev_valid0;
        valid_out <= prev_valid1;
        macroblock_out <= {row1, row2, row3, row4, row5, row6, row7, row8};
        row1 <= {block1, block2, block3, block4, block5, block6, block7, block8};
        row2 <= {block9, block10, block11, block12, block13, block14, block15, block16};
        row3 <= {block17, block18, block19, block20, block21, block22, block23, block24};
        row4 <= {block25, block26, block27, block28, block29, block30, block31, block32};
        row5 <= {block33, block34, block35, block36, block37, block38, block39, block40};
        row6 <= {block41, block42, block43, block44, block45, block46, block47, block48};
        row7 <= {block49, block50, block51, block52, block53, block54, block55, block56};
        row8 <= {block57, block58, block59, block60, block61, block62, block63, block64};
        if (rst) begin
            valid_out <= 0;
        end else if (valid_in) begin
            block1[0][0] <= {macroblock[0][0][23:16], macroblock[0][0][15:8], macroblock[0][0][7:0]};
            block1[0][1] <= {macroblock[0][1][23:16], macroblock[0][0][15:8], macroblock[0][0][7:0]};
            block1[1][0] <= {macroblock[1][0][23:16], macroblock[0][0][15:8], macroblock[0][0][7:0]};
            block1[1][1] <= {macroblock[1][1][23:16], macroblock[0][0][15:8], macroblock[0][0][7:0]};
            block2[0][0] <= {macroblock[0][2][23:16], macroblock[0][2][15:8], macroblock[0][2][7:0]};
            block2[0][1] <= {macroblock[0][3][23:16], macroblock[0][2][15:8], macroblock[0][2][7:0]};
            block2[1][0] <= {macroblock[1][2][23:16], macroblock[0][2][15:8], macroblock[0][2][7:0]};
            block2[1][1] <= {macroblock[1][3][23:16], macroblock[0][2][15:8], macroblock[0][2][7:0]};
            block3[0][0] <= {macroblock[0][4][23:16], macroblock[0][4][15:8], macroblock[0][4][7:0]};
            block3[0][1] <= {macroblock[0][5][23:16], macroblock[0][4][15:8], macroblock[0][4][7:0]};
            block3[1][0] <= {macroblock[1][4][23:16], macroblock[0][4][15:8], macroblock[0][4][7:0]};
            block3[1][1] <= {macroblock[1][5][23:16], macroblock[0][4][15:8], macroblock[0][4][7:0]};
            block4[0][0] <= {macroblock[0][6][23:16], macroblock[0][6][15:8], macroblock[0][6][7:0]};
            block4[0][1] <= {macroblock[0][7][23:16], macroblock[0][6][15:8], macroblock[0][6][7:0]};
            block4[1][0] <= {macroblock[1][6][23:16], macroblock[0][6][15:8], macroblock[0][6][7:0]};
            block4[1][1] <= {macroblock[1][7][23:16], macroblock[0][6][15:8], macroblock[0][6][7:0]};
            block5[0][0] <= {macroblock[0][8][23:16], macroblock[0][8][15:8], macroblock[0][8][7:0]};
            block5[0][1] <= {macroblock[0][9][23:16], macroblock[0][8][15:8], macroblock[0][8][7:0]};
            block5[1][0] <= {macroblock[1][8][23:16], macroblock[0][8][15:8], macroblock[0][8][7:0]};
            block5[1][1] <= {macroblock[1][9][23:16], macroblock[0][8][15:8], macroblock[0][8][7:0]};
            block6[0][0] <= {macroblock[0][10][23:16], macroblock[0][10][15:8], macroblock[0][10][7:0]};
            block6[0][1] <= {macroblock[0][11][23:16], macroblock[0][10][15:8], macroblock[0][10][7:0]};
            block6[1][0] <= {macroblock[1][10][23:16], macroblock[0][10][15:8], macroblock[0][10][7:0]};
            block6[1][1] <= {macroblock[1][11][23:16], macroblock[0][10][15:8], macroblock[0][10][7:0]};
            block7[0][0] <= {macroblock[0][12][23:16], macroblock[0][12][15:8], macroblock[0][12][7:0]};
            block7[0][1] <= {macroblock[0][13][23:16], macroblock[0][12][15:8], macroblock[0][12][7:0]};
            block7[1][0] <= {macroblock[1][12][23:16], macroblock[0][12][15:8], macroblock[0][12][7:0]};
            block7[1][1] <= {macroblock[1][13][23:16], macroblock[0][12][15:8], macroblock[0][12][7:0]};
            block8[0][0] <= {macroblock[0][14][23:16], macroblock[0][14][15:8], macroblock[0][14][7:0]};
            block8[0][1] <= {macroblock[0][15][23:16], macroblock[0][14][15:8], macroblock[0][14][7:0]};
            block8[1][0] <= {macroblock[1][14][23:16], macroblock[0][14][15:8], macroblock[0][14][7:0]};
            block8[1][1] <= {macroblock[1][15][23:16], macroblock[0][14][15:8], macroblock[0][14][7:0]};
            block9[0][0] <= {macroblock[2][0][23:16], macroblock[2][0][15:8], macroblock[2][0][7:0]};
            block9[0][1] <= {macroblock[2][1][23:16], macroblock[2][0][15:8], macroblock[2][0][7:0]};
            block9[1][0] <= {macroblock[3][0][23:16], macroblock[2][0][15:8], macroblock[2][0][7:0]};
            block9[1][1] <= {macroblock[3][1][23:16], macroblock[2][0][15:8], macroblock[2][0][7:0]};
            block10[0][0] <= {macroblock[2][2][23:16], macroblock[2][2][15:8], macroblock[2][2][7:0]};
            block10[0][1] <= {macroblock[2][3][23:16], macroblock[2][2][15:8], macroblock[2][2][7:0]};
            block10[1][0] <= {macroblock[3][2][23:16], macroblock[2][2][15:8], macroblock[2][2][7:0]};
            block10[1][1] <= {macroblock[3][3][23:16], macroblock[2][2][15:8], macroblock[2][2][7:0]};
            block11[0][0] <= {macroblock[2][4][23:16], macroblock[2][4][15:8], macroblock[2][4][7:0]};
            block11[0][1] <= {macroblock[2][5][23:16], macroblock[2][4][15:8], macroblock[2][4][7:0]};
            block11[1][0] <= {macroblock[3][4][23:16], macroblock[2][4][15:8], macroblock[2][4][7:0]};
            block11[1][1] <= {macroblock[3][5][23:16], macroblock[2][4][15:8], macroblock[2][4][7:0]};
            block12[0][0] <= {macroblock[2][6][23:16], macroblock[2][6][15:8], macroblock[2][6][7:0]};
            block12[0][1] <= {macroblock[2][7][23:16], macroblock[2][6][15:8], macroblock[2][6][7:0]};
            block12[1][0] <= {macroblock[3][6][23:16], macroblock[2][6][15:8], macroblock[2][6][7:0]};
            block12[1][1] <= {macroblock[3][7][23:16], macroblock[2][6][15:8], macroblock[2][6][7:0]};
            block13[0][0] <= {macroblock[2][8][23:16], macroblock[2][8][15:8], macroblock[2][8][7:0]};
            block13[0][1] <= {macroblock[2][9][23:16], macroblock[2][8][15:8], macroblock[2][8][7:0]};
            block13[1][0] <= {macroblock[3][8][23:16], macroblock[2][8][15:8], macroblock[2][8][7:0]};
            block13[1][1] <= {macroblock[3][9][23:16], macroblock[2][8][15:8], macroblock[2][8][7:0]};
            block14[0][0] <= {macroblock[2][10][23:16], macroblock[2][10][15:8], macroblock[2][10][7:0]};
            block14[0][1] <= {macroblock[2][11][23:16], macroblock[2][10][15:8], macroblock[2][10][7:0]};
            block14[1][0] <= {macroblock[3][10][23:16], macroblock[2][10][15:8], macroblock[2][10][7:0]};
            block14[1][1] <= {macroblock[3][11][23:16], macroblock[2][10][15:8], macroblock[2][10][7:0]};
            block15[0][0] <= {macroblock[2][12][23:16], macroblock[2][12][15:8], macroblock[2][12][7:0]};
            block15[0][1] <= {macroblock[2][13][23:16], macroblock[2][12][15:8], macroblock[2][12][7:0]};
            block15[1][0] <= {macroblock[3][12][23:16], macroblock[2][12][15:8], macroblock[2][12][7:0]};
            block15[1][1] <= {macroblock[3][13][23:16], macroblock[2][12][15:8], macroblock[2][12][7:0]};
            block16[0][0] <= {macroblock[2][14][23:16], macroblock[2][14][15:8], macroblock[2][14][7:0]};
            block16[0][1] <= {macroblock[2][15][23:16], macroblock[2][14][15:8], macroblock[2][14][7:0]};
            block16[1][0] <= {macroblock[3][14][23:16], macroblock[2][14][15:8], macroblock[2][14][7:0]};
            block16[1][1] <= {macroblock[3][15][23:16], macroblock[2][14][15:8], macroblock[2][14][7:0]};
            block17[0][0] <= {macroblock[4][0][23:16], macroblock[4][0][15:8], macroblock[4][0][7:0]};
            block17[0][1] <= {macroblock[4][1][23:16], macroblock[4][0][15:8], macroblock[4][0][7:0]};
            block17[1][0] <= {macroblock[5][0][23:16], macroblock[4][0][15:8], macroblock[4][0][7:0]};
            block17[1][1] <= {macroblock[5][1][23:16], macroblock[4][0][15:8], macroblock[4][0][7:0]};
            block18[0][0] <= {macroblock[4][2][23:16], macroblock[4][2][15:8], macroblock[4][2][7:0]};
            block18[0][1] <= {macroblock[4][3][23:16], macroblock[4][2][15:8], macroblock[4][2][7:0]};
            block18[1][0] <= {macroblock[5][2][23:16], macroblock[4][2][15:8], macroblock[4][2][7:0]};
            block18[1][1] <= {macroblock[5][3][23:16], macroblock[4][2][15:8], macroblock[4][2][7:0]};
            block19[0][0] <= {macroblock[4][4][23:16], macroblock[4][4][15:8], macroblock[4][4][7:0]};
            block19[0][1] <= {macroblock[4][5][23:16], macroblock[4][4][15:8], macroblock[4][4][7:0]};
            block19[1][0] <= {macroblock[5][4][23:16], macroblock[4][4][15:8], macroblock[4][4][7:0]};
            block19[1][1] <= {macroblock[5][5][23:16], macroblock[4][4][15:8], macroblock[4][4][7:0]};
            block20[0][0] <= {macroblock[4][6][23:16], macroblock[4][6][15:8], macroblock[4][6][7:0]};
            block20[0][1] <= {macroblock[4][7][23:16], macroblock[4][6][15:8], macroblock[4][6][7:0]};
            block20[1][0] <= {macroblock[5][6][23:16], macroblock[4][6][15:8], macroblock[4][6][7:0]};
            block20[1][1] <= {macroblock[5][7][23:16], macroblock[4][6][15:8], macroblock[4][6][7:0]};
            block21[0][0] <= {macroblock[4][8][23:16], macroblock[4][8][15:8], macroblock[4][8][7:0]};
            block21[0][1] <= {macroblock[4][9][23:16], macroblock[4][8][15:8], macroblock[4][8][7:0]};
            block21[1][0] <= {macroblock[5][8][23:16], macroblock[4][8][15:8], macroblock[4][8][7:0]};
            block21[1][1] <= {macroblock[5][9][23:16], macroblock[4][8][15:8], macroblock[4][8][7:0]};
            block22[0][0] <= {macroblock[4][10][23:16], macroblock[4][10][15:8], macroblock[4][10][7:0]};
            block22[0][1] <= {macroblock[4][11][23:16], macroblock[4][10][15:8], macroblock[4][10][7:0]};
            block22[1][0] <= {macroblock[5][10][23:16], macroblock[4][10][15:8], macroblock[4][10][7:0]};
            block22[1][1] <= {macroblock[5][11][23:16], macroblock[4][10][15:8], macroblock[4][10][7:0]};
            block23[0][0] <= {macroblock[4][12][23:16], macroblock[4][12][15:8], macroblock[4][12][7:0]};
            block23[0][1] <= {macroblock[4][13][23:16], macroblock[4][12][15:8], macroblock[4][12][7:0]};
            block23[1][0] <= {macroblock[5][12][23:16], macroblock[4][12][15:8], macroblock[4][12][7:0]};
            block23[1][1] <= {macroblock[5][13][23:16], macroblock[4][12][15:8], macroblock[4][12][7:0]};
            block24[0][0] <= {macroblock[4][14][23:16], macroblock[4][14][15:8], macroblock[4][14][7:0]};
            block24[0][1] <= {macroblock[4][15][23:16], macroblock[4][14][15:8], macroblock[4][14][7:0]};
            block24[1][0] <= {macroblock[5][14][23:16], macroblock[4][14][15:8], macroblock[4][14][7:0]};
            block24[1][1] <= {macroblock[5][15][23:16], macroblock[4][14][15:8], macroblock[4][14][7:0]};
            block25[0][0] <= {macroblock[6][0][23:16], macroblock[6][0][15:8], macroblock[6][0][7:0]};
            block25[0][1] <= {macroblock[6][1][23:16], macroblock[6][0][15:8], macroblock[6][0][7:0]};
            block25[1][0] <= {macroblock[7][0][23:16], macroblock[6][0][15:8], macroblock[6][0][7:0]};
            block25[1][1] <= {macroblock[7][1][23:16], macroblock[6][0][15:8], macroblock[6][0][7:0]};
            block26[0][0] <= {macroblock[6][2][23:16], macroblock[6][2][15:8], macroblock[6][2][7:0]};
            block26[0][1] <= {macroblock[6][3][23:16], macroblock[6][2][15:8], macroblock[6][2][7:0]};
            block26[1][0] <= {macroblock[7][2][23:16], macroblock[6][2][15:8], macroblock[6][2][7:0]};
            block26[1][1] <= {macroblock[7][3][23:16], macroblock[6][2][15:8], macroblock[6][2][7:0]};
            block27[0][0] <= {macroblock[6][4][23:16], macroblock[6][4][15:8], macroblock[6][4][7:0]};
            block27[0][1] <= {macroblock[6][5][23:16], macroblock[6][4][15:8], macroblock[6][4][7:0]};
            block27[1][0] <= {macroblock[7][4][23:16], macroblock[6][4][15:8], macroblock[6][4][7:0]};
            block27[1][1] <= {macroblock[7][5][23:16], macroblock[6][4][15:8], macroblock[6][4][7:0]};
            block28[0][0] <= {macroblock[6][6][23:16], macroblock[6][6][15:8], macroblock[6][6][7:0]};
            block28[0][1] <= {macroblock[6][7][23:16], macroblock[6][6][15:8], macroblock[6][6][7:0]};
            block28[1][0] <= {macroblock[7][6][23:16], macroblock[6][6][15:8], macroblock[6][6][7:0]};
            block28[1][1] <= {macroblock[7][7][23:16], macroblock[6][6][15:8], macroblock[6][6][7:0]};
            block29[0][0] <= {macroblock[6][8][23:16], macroblock[6][8][15:8], macroblock[6][8][7:0]};
            block29[0][1] <= {macroblock[6][9][23:16], macroblock[6][8][15:8], macroblock[6][8][7:0]};
            block29[1][0] <= {macroblock[7][8][23:16], macroblock[6][8][15:8], macroblock[6][8][7:0]};
            block29[1][1] <= {macroblock[7][9][23:16], macroblock[6][8][15:8], macroblock[6][8][7:0]};
            block30[0][0] <= {macroblock[6][10][23:16], macroblock[6][10][15:8], macroblock[6][10][7:0]};
            block30[0][1] <= {macroblock[6][11][23:16], macroblock[6][10][15:8], macroblock[6][10][7:0]};
            block30[1][0] <= {macroblock[7][10][23:16], macroblock[6][10][15:8], macroblock[6][10][7:0]};
            block30[1][1] <= {macroblock[7][11][23:16], macroblock[6][10][15:8], macroblock[6][10][7:0]};
            block31[0][0] <= {macroblock[6][12][23:16], macroblock[6][12][15:8], macroblock[6][12][7:0]};
            block31[0][1] <= {macroblock[6][13][23:16], macroblock[6][12][15:8], macroblock[6][12][7:0]};
            block31[1][0] <= {macroblock[7][12][23:16], macroblock[6][12][15:8], macroblock[6][12][7:0]};
            block31[1][1] <= {macroblock[7][13][23:16], macroblock[6][12][15:8], macroblock[6][12][7:0]};
            block32[0][0] <= {macroblock[6][14][23:16], macroblock[6][14][15:8], macroblock[6][14][7:0]};
            block32[0][1] <= {macroblock[6][15][23:16], macroblock[6][14][15:8], macroblock[6][14][7:0]};
            block32[1][0] <= {macroblock[7][14][23:16], macroblock[6][14][15:8], macroblock[6][14][7:0]};
            block32[1][1] <= {macroblock[7][15][23:16], macroblock[6][14][15:8], macroblock[6][14][7:0]};
            block33[0][0] <= {macroblock[8][0][23:16], macroblock[8][0][15:8], macroblock[8][0][7:0]};
            block33[0][1] <= {macroblock[8][1][23:16], macroblock[8][0][15:8], macroblock[8][0][7:0]};
            block33[1][0] <= {macroblock[9][0][23:16], macroblock[8][0][15:8], macroblock[8][0][7:0]};
            block33[1][1] <= {macroblock[9][1][23:16], macroblock[8][0][15:8], macroblock[8][0][7:0]};
            block34[0][0] <= {macroblock[8][2][23:16], macroblock[8][2][15:8], macroblock[8][2][7:0]};
            block34[0][1] <= {macroblock[8][3][23:16], macroblock[8][2][15:8], macroblock[8][2][7:0]};
            block34[1][0] <= {macroblock[9][2][23:16], macroblock[8][2][15:8], macroblock[8][2][7:0]};
            block34[1][1] <= {macroblock[9][3][23:16], macroblock[8][2][15:8], macroblock[8][2][7:0]};
            block35[0][0] <= {macroblock[8][4][23:16], macroblock[8][4][15:8], macroblock[8][4][7:0]};
            block35[0][1] <= {macroblock[8][5][23:16], macroblock[8][4][15:8], macroblock[8][4][7:0]};
            block35[1][0] <= {macroblock[9][4][23:16], macroblock[8][4][15:8], macroblock[8][4][7:0]};
            block35[1][1] <= {macroblock[9][5][23:16], macroblock[8][4][15:8], macroblock[8][4][7:0]};
            block36[0][0] <= {macroblock[8][6][23:16], macroblock[8][6][15:8], macroblock[8][6][7:0]};
            block36[0][1] <= {macroblock[8][7][23:16], macroblock[8][6][15:8], macroblock[8][6][7:0]};
            block36[1][0] <= {macroblock[9][6][23:16], macroblock[8][6][15:8], macroblock[8][6][7:0]};
            block36[1][1] <= {macroblock[9][7][23:16], macroblock[8][6][15:8], macroblock[8][6][7:0]};
            block37[0][0] <= {macroblock[8][8][23:16], macroblock[8][8][15:8], macroblock[8][8][7:0]};
            block37[0][1] <= {macroblock[8][9][23:16], macroblock[8][8][15:8], macroblock[8][8][7:0]};
            block37[1][0] <= {macroblock[9][8][23:16], macroblock[8][8][15:8], macroblock[8][8][7:0]};
            block37[1][1] <= {macroblock[9][9][23:16], macroblock[8][8][15:8], macroblock[8][8][7:0]};
            block38[0][0] <= {macroblock[8][10][23:16], macroblock[8][10][15:8], macroblock[8][10][7:0]};
            block38[0][1] <= {macroblock[8][11][23:16], macroblock[8][10][15:8], macroblock[8][10][7:0]};
            block38[1][0] <= {macroblock[9][10][23:16], macroblock[8][10][15:8], macroblock[8][10][7:0]};
            block38[1][1] <= {macroblock[9][11][23:16], macroblock[8][10][15:8], macroblock[8][10][7:0]};
            block39[0][0] <= {macroblock[8][12][23:16], macroblock[8][12][15:8], macroblock[8][12][7:0]};
            block39[0][1] <= {macroblock[8][13][23:16], macroblock[8][12][15:8], macroblock[8][12][7:0]};
            block39[1][0] <= {macroblock[9][12][23:16], macroblock[8][12][15:8], macroblock[8][12][7:0]};
            block39[1][1] <= {macroblock[9][13][23:16], macroblock[8][12][15:8], macroblock[8][12][7:0]};
            block40[0][0] <= {macroblock[8][14][23:16], macroblock[8][14][15:8], macroblock[8][14][7:0]};
            block40[0][1] <= {macroblock[8][15][23:16], macroblock[8][14][15:8], macroblock[8][14][7:0]};
            block40[1][0] <= {macroblock[9][14][23:16], macroblock[8][14][15:8], macroblock[8][14][7:0]};
            block40[1][1] <= {macroblock[9][15][23:16], macroblock[8][14][15:8], macroblock[8][14][7:0]};
            block41[0][0] <= {macroblock[10][0][23:16], macroblock[10][0][15:8], macroblock[10][0][7:0]};
            block41[0][1] <= {macroblock[10][1][23:16], macroblock[10][0][15:8], macroblock[10][0][7:0]};
            block41[1][0] <= {macroblock[11][0][23:16], macroblock[10][0][15:8], macroblock[10][0][7:0]};
            block41[1][1] <= {macroblock[11][1][23:16], macroblock[10][0][15:8], macroblock[10][0][7:0]};
            block42[0][0] <= {macroblock[10][2][23:16], macroblock[10][2][15:8], macroblock[10][2][7:0]};
            block42[0][1] <= {macroblock[10][3][23:16], macroblock[10][2][15:8], macroblock[10][2][7:0]};
            block42[1][0] <= {macroblock[11][2][23:16], macroblock[10][2][15:8], macroblock[10][2][7:0]};
            block42[1][1] <= {macroblock[11][3][23:16], macroblock[10][2][15:8], macroblock[10][2][7:0]};
            block43[0][0] <= {macroblock[10][4][23:16], macroblock[10][4][15:8], macroblock[10][4][7:0]};
            block43[0][1] <= {macroblock[10][5][23:16], macroblock[10][4][15:8], macroblock[10][4][7:0]};
            block43[1][0] <= {macroblock[11][4][23:16], macroblock[10][4][15:8], macroblock[10][4][7:0]};
            block43[1][1] <= {macroblock[11][5][23:16], macroblock[10][4][15:8], macroblock[10][4][7:0]};
            block44[0][0] <= {macroblock[10][6][23:16], macroblock[10][6][15:8], macroblock[10][6][7:0]};
            block44[0][1] <= {macroblock[10][7][23:16], macroblock[10][6][15:8], macroblock[10][6][7:0]};
            block44[1][0] <= {macroblock[11][6][23:16], macroblock[10][6][15:8], macroblock[10][6][7:0]};
            block44[1][1] <= {macroblock[11][7][23:16], macroblock[10][6][15:8], macroblock[10][6][7:0]};
            block45[0][0] <= {macroblock[10][8][23:16], macroblock[10][8][15:8], macroblock[10][8][7:0]};
            block45[0][1] <= {macroblock[10][9][23:16], macroblock[10][8][15:8], macroblock[10][8][7:0]};
            block45[1][0] <= {macroblock[11][8][23:16], macroblock[10][8][15:8], macroblock[10][8][7:0]};
            block45[1][1] <= {macroblock[11][9][23:16], macroblock[10][8][15:8], macroblock[10][8][7:0]};
            block46[0][0] <= {macroblock[10][10][23:16], macroblock[10][10][15:8], macroblock[10][10][7:0]};
            block46[0][1] <= {macroblock[10][11][23:16], macroblock[10][10][15:8], macroblock[10][10][7:0]};
            block46[1][0] <= {macroblock[11][10][23:16], macroblock[10][10][15:8], macroblock[10][10][7:0]};
            block46[1][1] <= {macroblock[11][11][23:16], macroblock[10][10][15:8], macroblock[10][10][7:0]};
            block47[0][0] <= {macroblock[10][12][23:16], macroblock[10][12][15:8], macroblock[10][12][7:0]};
            block47[0][1] <= {macroblock[10][13][23:16], macroblock[10][12][15:8], macroblock[10][12][7:0]};
            block47[1][0] <= {macroblock[11][12][23:16], macroblock[10][12][15:8], macroblock[10][12][7:0]};
            block47[1][1] <= {macroblock[11][13][23:16], macroblock[10][12][15:8], macroblock[10][12][7:0]};
            block48[0][0] <= {macroblock[10][14][23:16], macroblock[10][14][15:8], macroblock[10][14][7:0]};
            block48[0][1] <= {macroblock[10][15][23:16], macroblock[10][14][15:8], macroblock[10][14][7:0]};
            block48[1][0] <= {macroblock[11][14][23:16], macroblock[10][14][15:8], macroblock[10][14][7:0]};
            block48[1][1] <= {macroblock[11][15][23:16], macroblock[10][14][15:8], macroblock[10][14][7:0]};
            block49[0][0] <= {macroblock[12][0][23:16], macroblock[12][0][15:8], macroblock[12][0][7:0]};
            block49[0][1] <= {macroblock[12][1][23:16], macroblock[12][0][15:8], macroblock[12][0][7:0]};
            block49[1][0] <= {macroblock[13][0][23:16], macroblock[12][0][15:8], macroblock[12][0][7:0]};
            block49[1][1] <= {macroblock[13][1][23:16], macroblock[12][0][15:8], macroblock[12][0][7:0]};
            block50[0][0] <= {macroblock[12][2][23:16], macroblock[12][2][15:8], macroblock[12][2][7:0]};
            block50[0][1] <= {macroblock[12][3][23:16], macroblock[12][2][15:8], macroblock[12][2][7:0]};
            block50[1][0] <= {macroblock[13][2][23:16], macroblock[12][2][15:8], macroblock[12][2][7:0]};
            block50[1][1] <= {macroblock[13][3][23:16], macroblock[12][2][15:8], macroblock[12][2][7:0]};
            block51[0][0] <= {macroblock[12][4][23:16], macroblock[12][4][15:8], macroblock[12][4][7:0]};
            block51[0][1] <= {macroblock[12][5][23:16], macroblock[12][4][15:8], macroblock[12][4][7:0]};
            block51[1][0] <= {macroblock[13][4][23:16], macroblock[12][4][15:8], macroblock[12][4][7:0]};
            block51[1][1] <= {macroblock[13][5][23:16], macroblock[12][4][15:8], macroblock[12][4][7:0]};
            block52[0][0] <= {macroblock[12][6][23:16], macroblock[12][6][15:8], macroblock[12][6][7:0]};
            block52[0][1] <= {macroblock[12][7][23:16], macroblock[12][6][15:8], macroblock[12][6][7:0]};
            block52[1][0] <= {macroblock[13][6][23:16], macroblock[12][6][15:8], macroblock[12][6][7:0]};
            block52[1][1] <= {macroblock[13][7][23:16], macroblock[12][6][15:8], macroblock[12][6][7:0]};
            block53[0][0] <= {macroblock[12][8][23:16], macroblock[12][8][15:8], macroblock[12][8][7:0]};
            block53[0][1] <= {macroblock[12][9][23:16], macroblock[12][8][15:8], macroblock[12][8][7:0]};
            block53[1][0] <= {macroblock[13][8][23:16], macroblock[12][8][15:8], macroblock[12][8][7:0]};
            block53[1][1] <= {macroblock[13][9][23:16], macroblock[12][8][15:8], macroblock[12][8][7:0]};
            block54[0][0] <= {macroblock[12][10][23:16], macroblock[12][10][15:8], macroblock[12][10][7:0]};
            block54[0][1] <= {macroblock[12][11][23:16], macroblock[12][10][15:8], macroblock[12][10][7:0]};
            block54[1][0] <= {macroblock[13][10][23:16], macroblock[12][10][15:8], macroblock[12][10][7:0]};
            block54[1][1] <= {macroblock[13][11][23:16], macroblock[12][10][15:8], macroblock[12][10][7:0]};
            block55[0][0] <= {macroblock[12][12][23:16], macroblock[12][12][15:8], macroblock[12][12][7:0]};
            block55[0][1] <= {macroblock[12][13][23:16], macroblock[12][12][15:8], macroblock[12][12][7:0]};
            block55[1][0] <= {macroblock[13][12][23:16], macroblock[12][12][15:8], macroblock[12][12][7:0]};
            block55[1][1] <= {macroblock[13][13][23:16], macroblock[12][12][15:8], macroblock[12][12][7:0]};
            block56[0][0] <= {macroblock[12][14][23:16], macroblock[12][14][15:8], macroblock[12][14][7:0]};
            block56[0][1] <= {macroblock[12][15][23:16], macroblock[12][14][15:8], macroblock[12][14][7:0]};
            block56[1][0] <= {macroblock[13][14][23:16], macroblock[12][14][15:8], macroblock[12][14][7:0]};
            block56[1][1] <= {macroblock[13][15][23:16], macroblock[12][14][15:8], macroblock[12][14][7:0]};
            block57[0][0] <= {macroblock[14][0][23:16], macroblock[14][0][15:8], macroblock[14][0][7:0]};
            block57[0][1] <= {macroblock[14][1][23:16], macroblock[14][0][15:8], macroblock[14][0][7:0]};
            block57[1][0] <= {macroblock[15][0][23:16], macroblock[14][0][15:8], macroblock[14][0][7:0]};
            block57[1][1] <= {macroblock[15][1][23:16], macroblock[14][0][15:8], macroblock[14][0][7:0]};
            block58[0][0] <= {macroblock[14][2][23:16], macroblock[14][2][15:8], macroblock[14][2][7:0]};
            block58[0][1] <= {macroblock[14][3][23:16], macroblock[14][2][15:8], macroblock[14][2][7:0]};
            block58[1][0] <= {macroblock[15][2][23:16], macroblock[14][2][15:8], macroblock[14][2][7:0]};
            block58[1][1] <= {macroblock[15][3][23:16], macroblock[14][2][15:8], macroblock[14][2][7:0]};
            block59[0][0] <= {macroblock[14][4][23:16], macroblock[14][4][15:8], macroblock[14][4][7:0]};
            block59[0][1] <= {macroblock[14][5][23:16], macroblock[14][4][15:8], macroblock[14][4][7:0]};
            block59[1][0] <= {macroblock[15][4][23:16], macroblock[14][4][15:8], macroblock[14][4][7:0]};
            block59[1][1] <= {macroblock[15][5][23:16], macroblock[14][4][15:8], macroblock[14][4][7:0]};
            block60[0][0] <= {macroblock[14][6][23:16], macroblock[14][6][15:8], macroblock[14][6][7:0]};
            block60[0][1] <= {macroblock[14][7][23:16], macroblock[14][6][15:8], macroblock[14][6][7:0]};
            block60[1][0] <= {macroblock[15][6][23:16], macroblock[14][6][15:8], macroblock[14][6][7:0]};
            block60[1][1] <= {macroblock[15][7][23:16], macroblock[14][6][15:8], macroblock[14][6][7:0]};
            block61[0][0] <= {macroblock[14][8][23:16], macroblock[14][8][15:8], macroblock[14][8][7:0]};
            block61[0][1] <= {macroblock[14][9][23:16], macroblock[14][8][15:8], macroblock[14][8][7:0]};
            block61[1][0] <= {macroblock[15][8][23:16], macroblock[14][8][15:8], macroblock[14][8][7:0]};
            block61[1][1] <= {macroblock[15][9][23:16], macroblock[14][8][15:8], macroblock[14][8][7:0]};
            block62[0][0] <= {macroblock[14][10][23:16], macroblock[14][10][15:8], macroblock[14][10][7:0]};
            block62[0][1] <= {macroblock[14][11][23:16], macroblock[14][10][15:8], macroblock[14][10][7:0]};
            block62[1][0] <= {macroblock[15][10][23:16], macroblock[14][10][15:8], macroblock[14][10][7:0]};
            block62[1][1] <= {macroblock[15][11][23:16], macroblock[14][10][15:8], macroblock[14][10][7:0]};
            block63[0][0] <= {macroblock[14][12][23:16], macroblock[14][12][15:8], macroblock[14][12][7:0]};
            block63[0][1] <= {macroblock[14][13][23:16], macroblock[14][12][15:8], macroblock[14][12][7:0]};
            block63[1][0] <= {macroblock[15][12][23:16], macroblock[14][12][15:8], macroblock[14][12][7:0]};
            block63[1][1] <= {macroblock[15][13][23:16], macroblock[14][12][15:8], macroblock[14][12][7:0]};
            block64[0][0] <= {macroblock[14][14][23:16], macroblock[14][14][15:8], macroblock[14][14][7:0]};
            block64[0][1] <= {macroblock[14][15][23:16], macroblock[14][14][15:8], macroblock[14][14][7:0]};
            block64[1][0] <= {macroblock[15][14][23:16], macroblock[14][14][15:8], macroblock[14][14][7:0]};
            block64[1][1] <= {macroblock[15][15][23:16], macroblock[14][14][15:8], macroblock[14][14][7:0]};
        end
    end

endmodule
`default_nettype none
